library verilog;
use verilog.vl_types.all;
entity DUT2 is
end DUT2;
