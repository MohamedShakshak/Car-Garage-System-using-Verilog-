module car_garage(clk,reset,car_enter,car_out,car_count,garage_full,leds1,leds2,current_state,next_state);
  
  input clk,reset,car_enter,car_out;
  output  [5:0] car_count;
  output reg garage_full; // close 50 1  , Open < 50 0  
  output  [6:0]leds1,leds2;
 
  up_counter upCounter (clk,reset,car_enter,car_out,car_count); // Counter connection 
    
  parameter Max_cars=50; 
  
  parameter IDLE=2'b00,
            OPEN=2'b01,
            CLOSE=2'b10;
            
  output reg [1:0] current_state,next_state;
  
  
  always @(posedge clk or posedge reset)
  begin
    if(reset) begin
      current_state<=IDLE;
    end
  else
    current_state <= next_state;
  end 
  
  
 always @(*) 
 begin
   case(current_state)
     IDLE:begin
       if(car_enter) 
         next_state <=OPEN;
       else
         next_state=IDLE;
       end
       OPEN:begin
         if(car_enter && car_count < Max_cars)
           next_state=OPEN;
         else if(car_out)
           next_state=OPEN;
         else if(car_count == Max_cars)
           begin
             next_state=CLOSE;
         //    garage_full <=1'b1;
           end
	  else if(car_count == 6'b0)
		  next_state <= IDLE;
         end
         CLOSE:begin
           if(car_enter)
             begin
             next_state=CLOSE;
           // $display("GARAGE IS FULL ");
            end
           else if(car_out)
             begin
             /*  if(car_count == Max_cars )
                 begin
                   next_state <= CLOSE;
                   garage_full <= 1'b1;
                  // $display("GARAGE IS FULL ");
                 end*/              
             next_state=OPEN;
          //   garage_full <= 1'b0;
           end
         else if(reset)
           next_state=IDLE;
         end
           default: next_state = IDLE;
         endcase
       end  
       
       
        always @(posedge clk)
        begin
          case(current_state)
            IDLE: begin
              garage_full <=1'b0;
            end
            OPEN:begin
              garage_full <= 1'b0;
            end
            CLOSE : begin
              garage_full <= 1'b1;
              //$display("GARAGE IS FULL ");
            end
          endcase            
      end 
    // wire [6:0] led1,led2;
     counter_to_decoder CTD (clk,reset,car_count,leds1,leds2); 
   //  assign leds1=led1;
    // assign leds2=led2;
  
endmodule
