library verilog;
use verilog.vl_types.all;
entity DUT is
end DUT;
