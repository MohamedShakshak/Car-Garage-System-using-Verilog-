library verilog;
use verilog.vl_types.all;
entity up_counter_DUT is
end up_counter_DUT;
